LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.all;
USE IEEE.STD_LOGIC_UNSIGNED.all;

ENTITY RAM IS
PORT	(
	CLK		: IN	STD_LOGIC;
	RESET_NAI	: IN	STD_LOGIC;
	--
	RW_in		: IN	STD_LOGIC;
	DATA_in		: IN 	STD_LOGIC_VECTOR (7 DOWNTO 0);
	DATA_out	: OUT 	STD_LOGIC_VECTOR (7 DOWNTO 0);
	ADDRESS_in	: IN	STD_LOGIC_VECTOR (11 DOWNTO 0);
	RAM_SELECT_in	: IN	STD_LOGIC
	);
END RAM;

ARCHITECTURE TEST_RAM_ARCH OF RAM IS

SIGNAL	CLK_sig		: STD_LOGIC; 
SIGNAL	RESET_NAI_sig	: STD_LOGIC;
----
TYPE 	T_RAM IS ARRAY (0 TO 383) OF STD_LOGIC_VECTOR (7 DOWNTO 0);	
SIGNAL	RAM_DATA : T_RAM;
----
SIGNAL	DATA_in_sig		: STD_LOGIC_VECTOR (7 DOWNTO 0);
SIGNAL	DATA_out_sig		: STD_LOGIC_VECTOR (7 DOWNTO 0);
SIGNAL	ADDRESS_in_sig		: STD_LOGIC_VECTOR (11 DOWNTO 0);
SIGNAL	RW_in_sig		: STD_LOGIC;
SIGNAL	RAM_SELECT_in_sig	: STD_LOGIC;

BEGIN
DATA_in_sig		<= DATA_in;
DATA_out		<= DATA_out_sig;	
ADDRESS_in_sig		<= ADDRESS_in;
RW_in_sig		<= RW_in;
RAM_SELECT_in_sig	<= RAM_SELECT_in;

PROCESS(CLK,RESET_NAI)	
BEGIN
IF RESET_NAI = '0' THEN	
	DATA_out <= (OTHERS => '0');
ELSIF CLK'EVENT AND CLK = '1' THEN
	IF RAM_SELECT_in_sig = '1' THEN
		IF RW_in_sig = '0' THEN			-- write operation
			RAM_DATA (CONV_INTEGER(ADDRESS_in_sig)) <= DATA_in_sig;
		ELSIF RW_in_sig = '1' THEN		-- read operation
			DATA_out_sig <= RAM_DATA (CONV_INTEGER(ADDRESS_in_sig));
		END IF;	
	ELSIF RAM_SELECT_in_sig = '0' THEN 
		DATA_out_sig <= "ZZZZZZZZ";
	END IF;	
END IF;
END PROCESS;	

END TEST_RAM_ARCH;


